* SPICE3 file created from sawgen-fet-sky130.ext - technology: sky130A

.option scale=5000u

.subckt sawgen-fet-sky130 vdd Ri Rb vss Vd Vt Vb Csaw
X0 vss Vb vss sky130_fd_pr__res_high_po_0p35 l=1400
X1 Vb vdd vss sky130_fd_pr__res_high_po_0p35 l=1400
X2 vss Rb vss sky130_fd_pr__res_high_po_0p35 l=1400
X3 Csaw Ri vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=160
X4  Ri Ri vdd vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=3200 l=160
X5 Vd Vt Csaw vdd sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=3200 l=160
X6 Vt Vd vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=160
X7 Vd Vd vss vss sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=400 l=160
.ends
