**.subckt sawgen-bjt
C1 saw GND .1n m=1
Q1 saw vcur net2 2N3906 area=1 m=1
V1 VDD GND 10
R1 VDD vcur 1k m=1
R2 vcur GND 5k m=1
Q2 vt net1 GND 2N3904 area=1 m=1
Q3 net1 vt saw 2N3906 area=1 m=1
R3 vt GND 100 m=1
R4 VDD vt 100 m=1
R5 VDD net2 100k m=1
**** begin user architecture code


*
.model 2N3904 NPN(IS=1E-14 VAF=100   Bf=300 IKF=0.4 XTB=1.5 BR=4   CJC=4E-12  CJE=8E-12 RB=20 RC=0.1
+ RE=0.1   TR=250E-9  TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m mfg=Philips)

.model 2N3906 PNP(IS=1E-14 VAF=100   BF=200 IKF=0.4 XTB=1.5 BR=4   CJC=4.5E-12 CJE=10E-12 RB=20
+ RC=0.1 RE=0.1   TR=250E-9   TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40  Icrating=200m mfg=Philips)

.OPTION ABSTOL=1e-15.
.OPTION GMIN=1.0e-12.
.OPTION ITL1=1e5
.OPTION RSHUNT=1e12
.OPTION RELTOL=1e-5
.OPTION METHOD=gear
//.lib /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
//.include /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice


.ic V(saw)=0
.control
tran 1n 200u
plot V(saw) V(vcur) V(Vt)
.endc

**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
** flattened .save nodes
.end
