**.subckt sawgen-fet
V1 VDD GND 10
M1 vt vd GND 2N7002 m=1
M2 vd vt saw BSS84 m=1
R1 VDD vt 10k m=1
R2 vt GND 10k m=1
C2 saw GND 10n m=1
Q1 saw vcur net2 2N3906 area=1 m=1
R3 VDD vcur 1k m=1
R4 vcur GND 5k m=1
R7 net1 net2 1k m=1
Va net3 GND 0
Vb VDD net1 0
V2 GND VEE 10
M3 vd vd net3 2N7002 m=1
**** begin user architecture code


.model BSS84 VDMOS(pchan Rg=3 Vto=-2.1 Rd=2.4 Rs=1.8 Rb=3 Kp=.2 Cgdmax=.04n Cgdmin=.001n Cgs=.02n
+ Cjo=.01n Is=2p mfg=Philips Vds=-50 Ron=6000m Qg=1n)
.model 2N7002 VDMOS(Rg=3 Vto=1.6 Rd=0 Rs=.75 Rb=.14 Kp=.17 mtriode=1.25 Cgdmax=80p Cgdmin=12p
+ Cgs=50p Cjo=50p Is=.04p mfg=Fairchild Vds=60 Ron=2 Qg=1.5n)


.model 2N3904 NPN(IS=1E-14 VAF=100   Bf=300 IKF=0.4 XTB=1.5 BR=4   CJC=4E-12  CJE=8E-12 RB=20 RC=0.1
+ RE=0.1   TR=250E-9  TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m mfg=Philips)

.model 2N3906 PNP(IS=1E-14 VAF=100   BF=200 IKF=0.4 XTB=1.5 BR=4   CJC=4.5E-12 CJE=10E-12 RB=20
+ RC=0.1 RE=0.1   TR=250E-9   TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40  Icrating=200m mfg=Philips)

//.lib /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
//.include /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice


.ic V(saw)=0
.control
tran 1n 200u
plot V(saw) V(Vt) V(vd)
//plot V(vd)
//plot I(Vb)
.endc

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
.GLOBAL VEE
** flattened .save nodes
.end
