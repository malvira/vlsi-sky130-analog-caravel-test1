magic
tech sky130A
magscale 1 2
timestamp 1623526904
<< nwell >>
rect -338 -1897 338 1897
<< mvpmos >>
rect -80 -1600 80 1600
<< mvpdiff >>
rect -138 1588 -80 1600
rect -138 -1588 -126 1588
rect -92 -1588 -80 1588
rect -138 -1600 -80 -1588
rect 80 1588 138 1600
rect 80 -1588 92 1588
rect 126 -1588 138 1588
rect 80 -1600 138 -1588
<< mvpdiffc >>
rect -126 -1588 -92 1588
rect 92 -1588 126 1588
<< mvnsubdiff >>
rect -272 1819 272 1831
rect -272 1785 -164 1819
rect 164 1785 272 1819
rect -272 1773 272 1785
rect -272 1723 -214 1773
rect -272 -1723 -260 1723
rect -226 -1723 -214 1723
rect 214 1723 272 1773
rect -272 -1773 -214 -1723
rect 214 -1723 226 1723
rect 260 -1723 272 1723
rect 214 -1773 272 -1723
rect -272 -1785 272 -1773
rect -272 -1819 -164 -1785
rect 164 -1819 272 -1785
rect -272 -1831 272 -1819
<< mvnsubdiffcont >>
rect -164 1785 164 1819
rect -260 -1723 -226 1723
rect 226 -1723 260 1723
rect -164 -1819 164 -1785
<< poly >>
rect -80 1681 80 1697
rect -80 1647 -64 1681
rect 64 1647 80 1681
rect -80 1600 80 1647
rect -80 -1647 80 -1600
rect -80 -1681 -64 -1647
rect 64 -1681 80 -1647
rect -80 -1697 80 -1681
<< polycont >>
rect -64 1647 64 1681
rect -64 -1681 64 -1647
<< locali >>
rect -260 1785 -164 1819
rect 164 1785 260 1819
rect -260 1723 -226 1785
rect 226 1723 260 1785
rect -80 1647 -64 1681
rect 64 1647 80 1681
rect -126 1588 -92 1604
rect -126 -1604 -92 -1588
rect 92 1588 126 1604
rect 92 -1604 126 -1588
rect -80 -1681 -64 -1647
rect 64 -1681 80 -1647
rect -260 -1785 -226 -1723
rect 226 -1785 260 -1723
rect -260 -1819 -164 -1785
rect 164 -1819 260 -1785
<< viali >>
rect -64 1647 64 1681
rect -126 -1588 -92 1588
rect 92 -1588 126 1588
rect -64 -1681 64 -1647
<< metal1 >>
rect -76 1681 76 1687
rect -76 1647 -64 1681
rect 64 1647 76 1681
rect -76 1641 76 1647
rect -132 1588 -86 1600
rect -132 -1588 -126 1588
rect -92 -1588 -86 1588
rect -132 -1600 -86 -1588
rect 86 1588 132 1600
rect 86 -1588 92 1588
rect 126 -1588 132 1588
rect 86 -1600 132 -1588
rect -76 -1647 76 -1641
rect -76 -1681 -64 -1647
rect 64 -1681 76 -1647
rect -76 -1687 76 -1681
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -243 -1802 243 1802
string parameters w 16 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
