magic
tech sky130A
magscale 1 2
timestamp 1623535931
<< error_s >>
rect -626 2156 -620 2162
rect -540 2156 -534 2162
rect -2420 2150 -2414 2156
rect -632 2150 -626 2156
rect -534 2150 -528 2156
rect -2426 2144 -2420 2150
rect -2426 2070 -2420 2076
rect -2420 2064 -2414 2070
rect -632 2064 -626 2070
rect -534 2064 -528 2070
rect -626 2058 -620 2064
rect -540 2058 -534 2064
rect -1236 -90 -1220 -86
rect -1208 -118 -1192 -114
<< nwell >>
rect 80 3240 130 3310
<< locali >>
rect -2360 3560 -1940 3640
rect -430 3560 110 3640
rect -2410 -40 -2310 3160
rect -2116 3156 -2040 3160
rect -2130 -40 -2040 3156
rect -226 3042 -134 3158
rect 50 3050 130 3160
rect -620 1890 -540 2070
rect -1170 1830 -1110 1850
rect -618 1492 -544 1890
rect -1170 1170 -1110 1180
rect -130 -180 50 -90
<< viali >>
rect -620 2070 -540 2150
rect -1170 1850 -1110 1910
rect -1170 1180 -1110 1240
<< metal1 >>
rect -430 3560 130 3661
rect -417 3515 -343 3560
rect -419 3509 -341 3515
rect -419 3425 -341 3431
rect -2130 3280 -1079 3302
rect -2301 3200 -1079 3280
rect -2301 3199 -2158 3200
rect -2116 3199 -1079 3200
rect -2410 2150 -2310 3160
rect -2116 3156 -2040 3199
rect -2330 2070 -2310 2150
rect -2410 -40 -2310 2070
rect -2130 -40 -2040 3156
rect -1182 3059 -1079 3199
rect -1855 2850 -1785 2856
rect -1275 2850 -1205 3025
rect -200 3020 -130 3160
rect -1785 2780 -1205 2850
rect -1030 2848 -130 3020
rect -1855 2774 -1785 2780
rect -1275 2615 -1205 2780
rect -1036 2752 -130 2848
rect -1030 2610 -130 2752
rect -950 2600 -130 2610
rect -1679 2279 -1601 2285
rect -1679 2150 -1601 2201
rect -1679 2090 -1110 2150
rect -1679 270 -1601 2090
rect -1170 1916 -1110 2090
rect -632 2064 -626 2156
rect -534 2064 -528 2156
rect -1182 1910 -1098 1916
rect -1182 1850 -1170 1910
rect -1110 1850 -1098 1910
rect -1182 1844 -1098 1850
rect -1170 1246 -1110 1760
rect -1182 1240 -1098 1246
rect -1182 1180 -1170 1240
rect -1110 1180 -1098 1240
rect -1182 1174 -1098 1180
rect -1180 430 -1100 1100
rect -1210 350 -790 430
rect -710 350 -704 430
rect -1300 270 -1220 320
rect -1680 190 -1220 270
rect -1300 -90 -1220 190
rect -1040 280 -960 320
rect -1040 200 -360 280
rect -1040 -80 -960 200
rect -440 -90 -360 200
rect -200 -50 -130 2600
rect -90 430 -10 436
rect 20 430 100 3160
rect -10 350 100 430
rect -90 344 -10 350
rect 20 -40 100 350
rect -440 -170 50 -90
rect -1680 -340 -550 -220
<< via1 >>
rect -419 3431 -341 3509
rect -2420 2070 -2330 2150
rect -1855 2780 -1785 2850
rect -1679 2201 -1601 2279
rect -626 2150 -534 2156
rect -626 2070 -620 2150
rect -620 2070 -540 2150
rect -540 2070 -534 2150
rect -626 2064 -534 2070
rect -790 350 -710 430
rect -90 350 -10 430
<< metal2 >>
rect -1679 3431 -419 3509
rect -341 3431 -335 3509
rect -1861 2780 -1855 2850
rect -1785 2780 -1779 2850
rect -2420 2150 -2330 2156
rect -1855 2150 -1785 2780
rect -1679 2279 -1601 3431
rect -1685 2201 -1679 2279
rect -1601 2201 -1595 2279
rect -2330 2070 -626 2150
rect -2420 2064 -2330 2070
rect -790 430 -710 436
rect -710 350 -90 430
rect -10 350 -4 430
rect -790 344 -710 350
use sky130_fd_pr__pfet_g5v0d10v5_V4E25R  sky130_fd_pr__pfet_g5v0d10v5_V4E25R_0
timestamp 1623527015
transform 1 0 -1122 0 1 2817
box -338 -497 338 497
use sky130_fd_pr__diode_pd2nw_05v5_BQJJ87  sky130_fd_pr__diode_pd2nw_05v5_BQJJ87_0
timestamp 1623526904
transform 1 0 -1139 0 1 1721
box -321 -321 321 321
use sky130_fd_pr__diode_pd2nw_05v5_BQJJ87  sky130_fd_pr__diode_pd2nw_05v5_BQJJ87_1
timestamp 1623526904
transform 1 0 -1139 0 1 1061
box -321 -321 321 321
use sky130_fd_pr__nfet_g5v0d10v5_UQEUHA  sky130_fd_pr__nfet_g5v0d10v5_UQEUHA_0
timestamp 1623526904
transform 1 0 -1132 0 1 118
box -308 -458 308 458
use sky130_fd_pr__pfet_g5v0d10v5_TTPRW6  sky130_fd_pr__pfet_g5v0d10v5_TTPRW6_0
timestamp 1623526904
transform 1 0 -2222 0 1 1557
box -338 -1897 338 1897
use sky130_fd_pr__pfet_g5v0d10v5_TTPRW6  sky130_fd_pr__pfet_g5v0d10v5_TTPRW6_1
timestamp 1623526904
transform 1 0 -42 0 1 1557
box -338 -1897 338 1897
use sky130_fd_pr__res_high_po_0p35_QHYJR3  sky130_fd_pr__res_high_po_0p35_QHYJR3_0
timestamp 1623529677
transform 1 0 -1643 0 1 792
box -37 -1132 37 1132
use sky130_fd_pr__res_high_po_0p35_QHYJR3  sky130_fd_pr__res_high_po_0p35_QHYJR3_2
timestamp 1623529677
transform 0 -1 -1128 1 0 3597
box -37 -1132 37 1132
use sky130_fd_pr__res_high_po_0p35_QHYJR3  sky130_fd_pr__res_high_po_0p35_QHYJR3_1
timestamp 1623529677
transform 1 0 -583 0 1 792
box -37 -1132 37 1132
<< labels >>
flabel locali 80 3600 80 3600 1 FreeSans 480 0 0 0 VSS
port 1 n
flabel locali -2390 3130 -2390 3130 1 FreeSans 480 0 0 0 VDD
port 0 n
flabel locali 100 3100 100 3100 1 FreeSans 480 0 0 0 Vd
port 7 n
flabel locali -50 -160 -50 -160 1 FreeSans 480 0 0 0 Vt
port 5 n
flabel locali -210 3100 -210 3100 1 FreeSans 480 0 0 0 Csaw
port 4 n
flabel locali -2070 3120 -2070 3120 1 FreeSans 480 0 0 0 Ri
port 3 n
flabel locali -2330 3600 -2330 3600 1 FreeSans 480 0 0 0 Rb
port 2 n
flabel metal1 -1130 -320 -1130 -320 1 FreeSans 480 0 0 0 Vb
port 6 n
<< end >>
