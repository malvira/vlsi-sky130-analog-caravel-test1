magic
tech sky130A
timestamp 1606063140
<< nwell >>
rect -496 -248 496 248
<< mvpmos >>
rect -367 -100 -287 100
rect -258 -100 -178 100
rect -149 -100 -69 100
rect -40 -100 40 100
rect 69 -100 149 100
rect 178 -100 258 100
rect 287 -100 367 100
<< mvpdiff >>
rect -396 94 -367 100
rect -396 -94 -390 94
rect -373 -94 -367 94
rect -396 -100 -367 -94
rect -287 94 -258 100
rect -287 -94 -281 94
rect -264 -94 -258 94
rect -287 -100 -258 -94
rect -178 94 -149 100
rect -178 -94 -172 94
rect -155 -94 -149 94
rect -178 -100 -149 -94
rect -69 94 -40 100
rect -69 -94 -63 94
rect -46 -94 -40 94
rect -69 -100 -40 -94
rect 40 94 69 100
rect 40 -94 46 94
rect 63 -94 69 94
rect 40 -100 69 -94
rect 149 94 178 100
rect 149 -94 155 94
rect 172 -94 178 94
rect 149 -100 178 -94
rect 258 94 287 100
rect 258 -94 264 94
rect 281 -94 287 94
rect 258 -100 287 -94
rect 367 94 396 100
rect 367 -94 373 94
rect 390 -94 396 94
rect 367 -100 396 -94
<< mvpdiffc >>
rect -390 -94 -373 94
rect -281 -94 -264 94
rect -172 -94 -155 94
rect -63 -94 -46 94
rect 46 -94 63 94
rect 155 -94 172 94
rect 264 -94 281 94
rect 373 -94 390 94
<< mvnsubdiff >>
rect -463 209 463 215
rect -463 192 -409 209
rect 409 192 463 209
rect -463 186 463 192
rect -463 161 -434 186
rect -463 -161 -457 161
rect -440 -161 -434 161
rect 434 161 463 186
rect -463 -186 -434 -161
rect 434 -161 440 161
rect 457 -161 463 161
rect 434 -186 463 -161
rect -463 -192 463 -186
rect -463 -209 -409 -192
rect 409 -209 463 -192
rect -463 -215 463 -209
<< mvnsubdiffcont >>
rect -409 192 409 209
rect -457 -161 -440 161
rect 440 -161 457 161
rect -409 -209 409 -192
<< poly >>
rect -367 140 -287 148
rect -367 123 -359 140
rect -295 123 -287 140
rect -367 100 -287 123
rect -258 140 -178 148
rect -258 123 -250 140
rect -186 123 -178 140
rect -258 100 -178 123
rect -149 140 -69 148
rect -149 123 -141 140
rect -77 123 -69 140
rect -149 100 -69 123
rect -40 140 40 148
rect -40 123 -32 140
rect 32 123 40 140
rect -40 100 40 123
rect 69 140 149 148
rect 69 123 77 140
rect 141 123 149 140
rect 69 100 149 123
rect 178 140 258 148
rect 178 123 186 140
rect 250 123 258 140
rect 178 100 258 123
rect 287 140 367 148
rect 287 123 295 140
rect 359 123 367 140
rect 287 100 367 123
rect -367 -123 -287 -100
rect -367 -140 -359 -123
rect -295 -140 -287 -123
rect -367 -148 -287 -140
rect -258 -123 -178 -100
rect -258 -140 -250 -123
rect -186 -140 -178 -123
rect -258 -148 -178 -140
rect -149 -123 -69 -100
rect -149 -140 -141 -123
rect -77 -140 -69 -123
rect -149 -148 -69 -140
rect -40 -123 40 -100
rect -40 -140 -32 -123
rect 32 -140 40 -123
rect -40 -148 40 -140
rect 69 -123 149 -100
rect 69 -140 77 -123
rect 141 -140 149 -123
rect 69 -148 149 -140
rect 178 -123 258 -100
rect 178 -140 186 -123
rect 250 -140 258 -123
rect 178 -148 258 -140
rect 287 -123 367 -100
rect 287 -140 295 -123
rect 359 -140 367 -123
rect 287 -148 367 -140
<< polycont >>
rect -359 123 -295 140
rect -250 123 -186 140
rect -141 123 -77 140
rect -32 123 32 140
rect 77 123 141 140
rect 186 123 250 140
rect 295 123 359 140
rect -359 -140 -295 -123
rect -250 -140 -186 -123
rect -141 -140 -77 -123
rect -32 -140 32 -123
rect 77 -140 141 -123
rect 186 -140 250 -123
rect 295 -140 359 -123
<< locali >>
rect -457 192 -409 209
rect 409 192 457 209
rect 440 161 457 192
rect -367 123 -359 140
rect -295 123 -287 140
rect -258 123 -250 140
rect -186 123 -178 140
rect -149 123 -141 140
rect -77 123 -69 140
rect -40 123 -32 140
rect 32 123 40 140
rect 69 123 77 140
rect 141 123 149 140
rect 178 123 186 140
rect 250 123 258 140
rect 287 123 295 140
rect 359 123 367 140
rect -390 94 -373 102
rect -390 -102 -373 -94
rect -281 94 -264 102
rect -281 -102 -264 -94
rect -172 94 -155 102
rect -172 -102 -155 -94
rect -63 94 -46 102
rect -63 -102 -46 -94
rect 46 94 63 102
rect 46 -102 63 -94
rect 155 94 172 102
rect 155 -102 172 -94
rect 264 94 281 102
rect 264 -102 281 -94
rect 373 94 390 102
rect 373 -102 390 -94
rect -367 -140 -359 -123
rect -295 -140 -287 -123
rect -258 -140 -250 -123
rect -186 -140 -178 -123
rect -149 -140 -141 -123
rect -77 -140 -69 -123
rect -40 -140 -32 -123
rect 32 -140 40 -123
rect 69 -140 77 -123
rect 141 -140 149 -123
rect 178 -140 186 -123
rect 250 -140 258 -123
rect 287 -140 295 -123
rect 359 -140 367 -123
rect -457 -192 -440 -161
rect 440 -192 457 -161
rect -457 -209 -409 -192
rect 409 -209 457 -192
<< viali >>
rect -396 192 396 209
rect -457 161 -440 192
rect -457 19 -440 161
rect -359 123 -295 140
rect -250 123 -186 140
rect -141 123 -77 140
rect -32 123 32 140
rect 77 123 141 140
rect 186 123 250 140
rect 295 123 359 140
rect -390 10 -373 85
rect -281 -85 -264 -10
rect -172 10 -155 85
rect -63 -85 -46 -10
rect 46 10 63 85
rect 155 -85 172 -10
rect 264 10 281 85
rect 373 -85 390 -10
rect -359 -140 -295 -123
rect -250 -140 -186 -123
rect -141 -140 -77 -123
rect -32 -140 32 -123
rect 77 -140 141 -123
rect 186 -140 250 -123
rect 295 -140 359 -123
<< metal1 >>
rect -402 209 402 212
rect -460 192 -437 198
rect -460 19 -457 192
rect -440 19 -437 192
rect -402 192 -396 209
rect 396 192 402 209
rect -402 189 402 192
rect -365 140 -289 143
rect -365 123 -359 140
rect -295 123 -289 140
rect -365 120 -289 123
rect -256 140 -180 143
rect -256 123 -250 140
rect -186 123 -180 140
rect -256 120 -180 123
rect -147 140 -71 143
rect -147 123 -141 140
rect -77 123 -71 140
rect -147 120 -71 123
rect -38 140 38 143
rect -38 123 -32 140
rect 32 123 38 140
rect -38 120 38 123
rect 71 140 147 143
rect 71 123 77 140
rect 141 123 147 140
rect 71 120 147 123
rect 180 140 256 143
rect 180 123 186 140
rect 250 123 256 140
rect 180 120 256 123
rect 289 140 365 143
rect 289 123 295 140
rect 359 123 365 140
rect 289 120 365 123
rect -460 13 -437 19
rect -393 85 -370 91
rect -393 10 -390 85
rect -373 10 -370 85
rect -393 4 -370 10
rect -175 85 -152 91
rect -175 10 -172 85
rect -155 10 -152 85
rect -175 4 -152 10
rect 43 85 66 91
rect 43 10 46 85
rect 63 10 66 85
rect 43 4 66 10
rect 261 85 284 91
rect 261 10 264 85
rect 281 10 284 85
rect 261 4 284 10
rect -284 -10 -261 -4
rect -284 -85 -281 -10
rect -264 -85 -261 -10
rect -284 -91 -261 -85
rect -66 -10 -43 -4
rect -66 -85 -63 -10
rect -46 -85 -43 -10
rect -66 -91 -43 -85
rect 152 -10 175 -4
rect 152 -85 155 -10
rect 172 -85 175 -10
rect 152 -91 175 -85
rect 370 -10 393 -4
rect 370 -85 373 -10
rect 390 -85 393 -10
rect 370 -91 393 -85
rect -365 -123 -289 -120
rect -365 -140 -359 -123
rect -295 -140 -289 -123
rect -365 -143 -289 -140
rect -256 -123 -180 -120
rect -256 -140 -250 -123
rect -186 -140 -180 -123
rect -256 -143 -180 -140
rect -147 -123 -71 -120
rect -147 -140 -141 -123
rect -77 -140 -71 -123
rect -147 -143 -71 -140
rect -38 -123 38 -120
rect -38 -140 -32 -123
rect 32 -140 38 -123
rect -38 -143 38 -140
rect 71 -123 147 -120
rect 71 -140 77 -123
rect 141 -140 147 -123
rect 71 -143 147 -140
rect 180 -123 256 -120
rect 180 -140 186 -123
rect 250 -140 256 -123
rect 180 -143 256 -140
rect 289 -123 365 -120
rect 289 -140 295 -123
rect 359 -140 365 -123
rect 289 -143 365 -140
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -448 -201 448 201
string parameters w 2.00 l 0.80 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl -45 viagr 0 viagt 90 viagb 0 viagate 100 viadrn -40 viasrc +40
string library sky130
<< end >>
