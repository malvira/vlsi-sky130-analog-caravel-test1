**.subckt sawgen-fet-sky130_tb
V1 VDD GND 10
x1 VDD cur cur GND Vd Vt Vt saw sawgen-fet-sky130
C1 saw GND 1n m=1
**** begin user architecture code


.model BSS84 VDMOS(pchan Rg=3 Vto=-2.1 Rd=2.4 Rs=1.8 Rb=3 Kp=.2 Cgdmax=.04n Cgdmin=.001n Cgs=.02n
+ Cjo=.01n Is=2p mfg=Philips Vds=-50 Ron=6000m Qg=1n)
.model 2N7002 VDMOS(Rg=3 Vto=1.6 Rd=0 Rs=.75 Rb=.14 Kp=.17 mtriode=1.25 Cgdmax=80p Cgdmin=12p
+ Cgs=50p Cjo=50p Is=.04p mfg=Fairchild Vds=60 Ron=2 Qg=1.5n)


.model 2N3904 NPN(IS=1E-14 VAF=100   Bf=300 IKF=0.4 XTB=1.5 BR=4   CJC=4E-12  CJE=8E-12 RB=20 RC=0.1
+ RE=0.1   TR=250E-9  TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40 Icrating=200m mfg=Philips)

.model 2N3906 PNP(IS=1E-14 VAF=100   BF=200 IKF=0.4 XTB=1.5 BR=4   CJC=4.5E-12 CJE=10E-12 RB=20
+ RC=0.1 RE=0.1   TR=250E-9   TF=350E-12 ITF=1 VTF=2 XTF=3 Vceo=40  Icrating=200m mfg=Philips)

//.include /usr/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_g5v0d10v5.pm3.spice
//.include /usr/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__res_high_po_0p35.model.spice

.lib /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice


.ic V(saw)=0
.control
tran 10n 200u
plot V(saw) V(cur) V(vt) V(vd)
//V(Vt) V(vd)
//plot V(vd)
//plot I(Vb)
.endc

**** end user architecture code
**.ends

* expanding   symbol:  sawgen-fet-sky130.sym # of pins=8
* sym_path:
*+ /home/malvira/repos/asic/projects/vlsi-sky130-analog-caravel-test1/xschem/sawgen-fet-sky130.sym
* sch_path:
*+ /home/malvira/repos/asic/projects/vlsi-sky130-analog-caravel-test1/xschem/sawgen-fet-sky130.sch
.subckt sawgen-fet-sky130  vdd Ri Rb vss Vd vt vb Csaw
*.ipin VDD
*.ipin VSS
*.iopin cur
*.iopin VSS
*.iopin Rb
*.iopin Ri
*.iopin Csaw
*.iopin Vt
*.iopin Vb
*.iopin Vd
XM5 Ri Ri VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 Csaw Ri VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XR8 VSS Rb VSS sky130_fd_pr__res_high_po_0p35 W=0.35 L=20 mult=1 m=1
XM1 Vd Vt Csaw VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=16 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 Vt Vd VSS GND sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XR3 Vb VDD VSS sky130_fd_pr__res_high_po_0p35 W=0.35 L=20 mult=1 m=1
XR4 VSS Vb VSS sky130_fd_pr__res_high_po_0p35 W=0.35 L=20 mult=1 m=1
D1 Vd net1 sky130_fd_pr__diode_pw2nd_05v5 area=1
D2 net1 VSS sky130_fd_pr__diode_pw2nd_05v5 area=1
.ends

.GLOBAL VDD
.GLOBAL GND
** flattened .save nodes
.end
